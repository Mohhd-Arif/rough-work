0,1
date,1568698184067
totalApiHit,1
totalLocHit,1
fetchLocHit,1
updateLocHit,0
trackerList,"{""shjckhww"":1}"
